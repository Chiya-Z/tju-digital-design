module mod_pos (
	input 	a, b, c, d,
	output	out1, out2
);

	// 代码量预计1行
	mod_a DUT(a, b, c, d, out1, out2);

endmodule
