module notgate (
	input 	in,    
	output 	out	
);

	// 代码量预计1行
	assign out = ~in;

endmodule
