module Kmap1(
    input   a,
    input   b,
    input   c,
    output  out
);

	// 代码量预计1行
    assign out = (a | b | c);

endmodule
