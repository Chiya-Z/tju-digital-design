module wire4 (
	input 	a, b, c,    
	output 	w, x, y, z	
);

	// 代码量预计4行
	assign w = a;
	assign x = b;
	assign y = b;
	assign z = c;

endmodule
