module wire1 (
	input 	in,    
	output 	out	
);

	// 代码量预计1行
	assign out = in;

endmodule