module compare (
	input 	[7 : 0] a, b,
	output	[2 : 0] flag, flag_s
);

	// 代码量预计3行
	assign {flag[0], flag_s[0]} = {2{(a == b)}};
	assign {flag[2], flag[1]} = (a < b)? 2'b01 : ((a > b)? 2'b10 : 2'b00);
	assign {flag_s[2], flag_s[1]} = ({a[0], b[0]} == 2'b10)? 2'b01 : 
									 (({a[0], b[0]} == 2'b01)? 2'b10 : (({a[0], b[0]} == 2'b00 && (a[6:0] < b[6:0]))? 2'b01 : (({a[0], b[0]} == 2'b00 && (a[6:0] > b[6:0]))? 2'b10 : (({a[0], b[0]} == 2'b11 && (a[6:0] > b[6:0]))? 2'b01 : (({a[0], b[0]} == 2'b11 && (a[6:0] < b[6:0]))? 2'b10 : 2'b00)))));
									

endmodule
