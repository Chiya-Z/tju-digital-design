module mod_name (
	input 	a, b, c, d,
	output	out1, out2
);

	// 代码量预计1行
	mod_a DUT(.a(a), .b(b), .c(c), .d(d), .out1(out1), .out2(out2));

endmodule
