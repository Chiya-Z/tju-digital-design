module andgate (
	input 	a,
	input	b,    
	output 	out	
);

	// 代码量预计1行
	assign out = a & b;

endmodule
