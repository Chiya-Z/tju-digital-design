module vector_concat (
	input 	[4 : 0] a, b, c, d, e, f,
	output	[7 : 0]	w, x, y, z
);

	// 代码量预计1行
	assign { w, x, y, z } = { a, b, c, d, e, f, 2'b11 };

endmodule
