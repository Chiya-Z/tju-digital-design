module vector_gate (
	input 	[2 : 0] a, b,
	output	[2 : 0] out_or_bitwise,
	output			out_or_logical,
	output	[5 : 0] out_not
);

	// 代码量预计3行
	assign out_or_bitwise = a | b;
    assign out_or_logical = a || b;
    assign out_not = {~b, ~a};

endmodule
